// Inspired by https://kastner.ucsd.edu/wp-content/uploads/2023/01/admin/isfpga23-turnon.pdf.
// See Figure 3.


